/* ****************************************************************************
 * Copyright(c) 2011-2016, Intel Corporation
 *
 * Redistribution and use in source and binary forms, with or without
 * modification, are permitted provided that the following conditions are met:
 *
 * * Redistributions of source code must retain the above copyright notice,
 * this list of conditions and the following disclaimer.
 * * Redistributions in binary form must reproduce the above copyright notice,
 * this list of conditions and the following disclaimer in the documentation
 * and/or other materials provided with the distribution.
 * * Neither the name of Intel Corporation nor the names of its contributors
 * may be used to endorse or promote products derived from this software
 * without specific prior written permission.
 *
 * THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
 * AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
 * IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
 * ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT OWNER OR CONTRIBUTORS BE
 * LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
 * CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
 * SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
 * INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
 * CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
 * ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
 * POSSIBILITY OF SUCH DAMAGE.
 *
 * **************************************************************************
 *
 * Module Info: CCI Transactions Logger
 * Language   : System{Verilog}
 * Owner      : Rahul R Sharma
 *              rahul.r.sharma@intel.com
 *              Intel Corporation
 *
 */

import ase_pkg::*;
import ccip_if_pkg::*;

`include "platform.vh"

module ccip_logger
  #(
    parameter LOGNAME   = "CHANGE_MY_NAME.log"
    )
   (
    // Configure enable
    input logic finish_logger,
    // Buffer message injection
    input logic log_timestamp_en,
    input logic log_string_en,
    ref string 	log_string,
    //////////////////////////////////////////////////////////
    // CCI interface
    input logic clk,
    input logic SoftReset,
    input 	t_if_ccip_Rx ccip_rx,
    input 	t_if_ccip_Tx ccip_tx
    );

   
   /*
    * ASE Hardware Interface (CCI) logger
    * - Logs CCI transaction into a transactions.tsv file
    * - Watch for "*valid", and write transaction to log name
    */
   // Log file descriptor
   int 					    log_fd;

   // Reset management
   logic 				    SoftReset_q;

   // Registers for comparing previous states
   always @(posedge clk) begin
      SoftReset_q	<= SoftReset;
   end

   // Config header
   t_ccip_c0_ReqMmioHdr C0RxMmioHdr;
   assign C0RxMmioHdr = t_ccip_c0_ReqMmioHdr'(ccip_rx.c0.hdr);

   // Umsg header
   UMsgHdr_t C0RxUMsgHdr;
   assign C0RxUMsgHdr = UMsgHdr_t'(ccip_rx.c0.hdr);

   
   /*
    * Buffer channels, request and response types
    */
   // Print Channel function
   function string print_channel (t_ccip_vc vc_sel);
      begin
   	 case (vc_sel)
   	   eVC_VA  : return "VA ";
   	   eVC_VL0 : return "VL0";
   	   eVC_VH0 : return "VH0";
   	   eVC_VH1 : return "VH1";
   	 endcase
      end
   endfunction

   // Print Req Type - CH0
   function string print_c0_reqtype (t_ccip_c0_ReqMemHdr req);
      begin
	 case (req)
	   eREQ_RDLINE_S   : return "Rd_S       ";
	   eREQ_RDLINE_I   : return "Rd_I       ";
	   default        : return "** ERROR %m : eREQ-CH0 unindentified **" ;
	 endcase
      end
   endfunction
   
   // Print req type - CH1
   function string print_c1_reqtype (t_ccip_c1_ReqMemHdr req);
      begin
	 case (req)
	   eREQ_WRLINE_I   : return "Wr_I       ";
	   eREQ_WRLINE_M   : return "Wr_M       ";
	   eREQ_WRFENCE    : return "WrFence    ";
	   eREQ_INTR       : return "IntrReq    ";
	   default         : return "** ERROR %m : eREQ-CH1 unindentified **" ;
	 endcase
      end
   endfunction

   // Print CH0 response type
   function string print_c0_resptype (t_ccip_c0_rsp resp);
      begin
	 case (resp)
	   eRSP_RDLINE     : return "RdResp     ";
	   default         : return "** ERROR %m : eRSP-CH0 unindentified **" ;
	 endcase
      end
   endfunction

   // Print CH1 response type
   function string print_c1_resptype (t_ccip_c1_rsp resp);
      begin
	 case (resp)
	   eRSP_WRLINE     : return "WrResp     ";
	   eRSP_WRFENCE    : return "WrFenceResp";
	   eRSP_INTR       : return "IntrResp   ";
	   default         : return "** ERROR %m : eRSP-CH1 unindentified **" ;
	 endcase
      end
   endfunction

   
   // Print CL number (in Request)
   function string print_cllen (t_ccip_clLen len);
      begin
	 case (len)
	   eCL_LEN_1 : return "#1CL";
	   eCL_LEN_2 : return "#2CL";
	   eCL_LEN_4 : return "#4CL";
	   default : return "** ERROR %m : clLen unindentified **" ;
	 endcase
      end
   endfunction

   
   // Print CL number (in Response)
   function string print_clnum (t_ccip_clNum num);
      begin
	 case (num)
	   2'b00 : return "#1CL";
	   2'b01 : return "#2CL";
	   2'b10 : return "#3CL";
	   2'b11 : return "#4CL";
	 endcase
      end
   endfunction

   
   // Print CSR data
   function string csr_data(int num_bytes, logic [CCIP_DATA_WIDTH-1:0] rx0_data);
      string str_4;
      string str_8;
      string str_64;
      begin
	 case (num_bytes)
	   4 :
	     begin
		str_4.hextoa(rx0_data[31:0]);
		return str_4;
	     end
	   8 :
	     begin
		str_8.hextoa(rx0_data[63:0]);
		return str_8;
	     end
	   64 :
	     begin
		str_64.hextoa(rx0_data[511:0]);
		return str_64;
	     end
	 endcase
      end
   endfunction

   
   // MMIO Request length
   function int mmioreq_length (logic [1:0] mmio_len);
      begin
	 case (mmio_len)
	   2'b00 : return 4;
	   2'b01 : return 8;
	   2'b10 : return 64;
	 endcase
      end
   endfunction // mmioreq_length

   
   // Space generator - formatting help
   function string ret_spaces (int num);
      string spaces;
      int    ii;
      begin
	 spaces = "";
	 for (ii = 0; ii < num; ii = ii + 1) begin
	    spaces = {spaces, " "};
	 end
	 return spaces;
      end
   endfunction


   /*
    * Function checks 
    */ 
   // Is a Read Request
   function logic isRdLineRequest(t_ccip_c0_req req);
      begin
	 if ((req == eREQ_RDLINE_I)||(req == eREQ_RDLINE_S)) 
	   return 1;
	 else
	   return 0;
      end
   endfunction
   
   // Is a Write Request
   function logic isWrLineRequest(t_ccip_c1_req req);
      begin
	 if ((req == eREQ_WRLINE_I)||(req == eREQ_WRLINE_M)) 
	   return 1;
	 else
	   return 0;
      end
   endfunction

   // Is a Write Fence Request
   function logic isWrFenceRequest(t_ccip_c1_req req);
      begin
	 if (req == eREQ_WRFENCE)
	   return 1;
	 else
	   return 0;
      end
   endfunction

   // Is a Intr Request
   function logic isIntrRequest(t_ccip_c1_req req);
      begin
	 if (req == eREQ_INTR)
	   return 1;
	 else
	   return 0;
      end
   endfunction
   
   // Is a Read Response
   function logic isRdLineResponse(t_ccip_c0_rsp rsp);
      begin
	 if (rsp == eRSP_RDLINE)
	   return 1;
	 else
	   return 0;
      end
   endfunction
   
   // Is a Umsg Response
   function logic isUmsgResponse(t_ccip_c0_rsp rsp);
      begin
	 if (rsp == eRSP_UMSG)
	   return 1;
	 else
	   return 0;
      end
   endfunction
   
   // Is a Write Response
   function logic isWrLineResponse(t_ccip_c1_rsp rsp);
      begin
	 if (rsp == eRSP_WRLINE)
	   return 1;
	 else
	   return 0;
      end
   endfunction
   
   // Is a Write Fence Response
   function logic isWrFenceResponse(t_ccip_c1_rsp rsp);
      begin
	 if (rsp == eRSP_WRFENCE)
	   return 1;
	 else
	   return 0;
      end
   endfunction
   

   /*
    * Watcher process
    */
   initial begin : logger_proc
      // Display
      $display("SIM-SV: Transaction Logger started");

      // Open transactions.tsv file
      log_fd = $fopen(LOGNAME, "w");

      // Watch CCI port
      forever begin
	 // Indicate Software controlled reset
	 if (SoftReset_q != SoftReset) begin
	    if (cfg.enable_cl_view) begin
	       $display("%d\tSoftReset toggled from %b to %b\n", $time, SoftReset_q, SoftReset);
	    end
	    $fwrite(log_fd, "%d\tSoftReset toggled from %b to %b\n", $time, SoftReset_q, SoftReset);
	 end
	 // Buffer messages
	 if (log_string_en) begin
	    if (log_timestamp_en) begin
	       $fwrite(log_fd, "-----------------------------------------------------\n");
	       $fwrite(log_fd, "%d\t%s\n", $time, log_string);
	    end
	    else begin
	       $fwrite(log_fd, "-----------------------------------------------------\n");
	       $fwrite(log_fd, "%s\n", log_string);	       
	    end
	 end
	 /////////////////////// CONFIG CHANNEL TRANSACTIONS //////////////////////////
	 /******************* MMIO Write Request *******************/
	 if (ccip_rx.c0.mmioWrValid) begin
	    if (cfg.enable_cl_view)  $display("%d\t   \tMMIOWrReq   \t%x\t%d bytes\t%s\n",
					      $time,
					      C0RxMmioHdr.address,
					      mmioreq_length(C0RxMmioHdr.length),
					      csr_data(mmioreq_length(C0RxMmioHdr.length), ccip_rx.c0.data)  );
	    $fwrite(log_fd, "%d\t   \tMMIOWrReq   \t  \t%x\t%d bytes\t%s\n",
					      $time,
					      C0RxMmioHdr.address,
					      mmioreq_length(C0RxMmioHdr.length),
					      csr_data(mmioreq_length(C0RxMmioHdr.length), ccip_rx.c0.data)  );
	 end
	 /******************* MMIO Read Request *******************/
	 if (ccip_rx.c0.mmioRdValid) begin
	    if (cfg.enable_cl_view) $display("%d\t   \tMMIORdReq   \t%x\t%x\t%d bytes\n",
	    				     $time,
	    				     C0RxMmioHdr.tid,
	    				     C0RxMmioHdr.address,
	    				     mmioreq_length(C0RxMmioHdr.length));
	    $fwrite(log_fd, "%d\t   \tMMIORdReq   \t%x\t%x\t%d bytes\n",
	    	    $time,
	    	    C0RxMmioHdr.tid,
	    	    C0RxMmioHdr.address,
	    	    mmioreq_length(C0RxMmioHdr.length));
	 end
	 //////////////////////// C0 TX CHANNEL TRANSACTIONS //////////////////////////
	 /******************* AFU -> MEM Read Request *****************/
	 if (ccip_tx.c0.valid && isRdLineRequest(ccip_tx.c0.hdr.req_type) ) begin
	    if (cfg.enable_cl_view) $display("%d\t%s\t%s\t%x\t%x\t%s",
	 				     $time,
	 				     print_channel(ccip_tx.c0.hdr.vc_sel),
	 				     print_c0_reqtype(ccip_tx.c0.hdr.req_type),
	 				     ccip_tx.c0.hdr.mdata,
	 				     ccip_tx.c0.hdr.address,
					     print_cllen(ccip_tx.c0.hdr.cl_len));
	    $fwrite(log_fd, "%d\t%s\t%s\t%x\t%x\t%s\n",
	 				     $time,
	 				     print_channel(ccip_tx.c0.hdr.vc_sel),
	 				     print_c0_reqtype(ccip_tx.c0.hdr.req_type),
	 				     ccip_tx.c0.hdr.mdata,
	 				     ccip_tx.c0.hdr.address,
					     print_cllen(ccip_tx.c0.hdr.cl_len));
	 end
	 //////////////////////// C1 TX CHANNEL TRANSACTIONS //////////////////////////
	 /******************* AFU -> MEM Write Request *****************/
	 if (ccip_tx.c1.valid && isWrLineRequest(ccip_tx.c1.hdr.req_type)) begin
	    if (cfg.enable_cl_view) $display("%d\t%s\t%s\t%x\t%x\t%x\t%s",
	 				     $time,
	 				     print_channel(ccip_tx.c1.hdr.vc_sel),
	 				     print_c1_reqtype(ccip_tx.c1.hdr.req_type),
	 				     ccip_tx.c1.hdr.mdata,
	 				     ccip_tx.c1.hdr.address,
	 				     ccip_tx.c1.data,
					     print_clnum(ccip_tx.c1.hdr.cl_len));
	    $fwrite(log_fd, "%d\t%s\t%s\t%x\t%x\t%x\t%s\n",
	 				     $time,
	 				     print_channel(ccip_tx.c1.hdr.vc_sel),
	 				     print_c1_reqtype(ccip_tx.c1.hdr.req_type),
	 				     ccip_tx.c1.hdr.mdata,
	 				     ccip_tx.c1.hdr.address,
	 				     ccip_tx.c1.data,
					     print_clnum(ccip_tx.c1.hdr.cl_len));
	 end // if (ccip_tx.c1.valid && (ccip_tx.c1.hdr.req_type != eREQ_WRFENCE))
	 if (ccip_tx.c1.valid && isWrFenceRequest(ccip_tx.c1.hdr.req_type)) begin
	    if (cfg.enable_cl_view) $display("%d\t%s\tWrFence \t%x\n",
					     $time,
					     print_channel(ccip_tx.c1.hdr.vc_sel),
					     ccip_tx.c1.hdr.mdata);
	    $fwrite(log_fd, "%d\t%s\tWrFence \t%x\n",
		    $time,
		    print_channel(ccip_tx.c1.hdr.vc_sel),
		    ccip_tx.c1.hdr.mdata);
	 end	 
	 //////////////////////// C2 TX CHANNEL TRANSACTIONS //////////////////////////
	 /********************** MMIO Read Response ********************/
	 if (ccip_tx.c2.mmioRdValid) begin
	    if (cfg.enable_cl_view) $display("%d\t   \tMMIORdRsp   \t%x\t%x\n",
					     $time,
					     ccip_tx.c2.hdr.tid,
					     ccip_tx.c2.data);
	    $fwrite(log_fd, "%d\t   \tMMIORdRsp   \t%x\t%x\n",
		    $time,
		    ccip_tx.c2.hdr.tid,
		    ccip_tx.c2.data);
	 end
	 //////////////////////// C0 RX CHANNEL TRANSACTIONS //////////////////////////
	 /******************* MEM -> AFU Read Response *****************/
	 if (ccip_rx.c0.rspValid && isRdLineResponse(ccip_rx.c0.hdr.resp_type)) begin
	    if (cfg.enable_cl_view) $display("%d\t%s\t%s\t%x\t%s\t%x",
	 				     $time,
	 				     print_channel(ccip_rx.c0.hdr.vc_used),
	 				     print_c0_resptype(ccip_rx.c0.hdr.resp_type),
	 				     ccip_rx.c0.hdr.mdata,
					     print_clnum(ccip_rx.c0.hdr.cl_num),
	 				     ccip_rx.c0.data);
	    $fwrite(log_fd, "%d\t%s\t%s\t%x\t%s\t%x\n",
	 				     $time,
	 				     print_channel(ccip_rx.c0.hdr.vc_used),
	 				     print_c0_resptype(ccip_rx.c0.hdr.resp_type),
	 				     ccip_rx.c0.hdr.mdata,
					     print_clnum(ccip_rx.c0.hdr.cl_num),
	 				     ccip_rx.c0.data);
	 end // if (ccip_tx.c0.rspValid && (ccip_rx.c0.hdr.resptype == eRSP_RDLINE)) 
	 /*************** SW -> MEM -> AFU Unordered Message  *************/
	 if (ccip_rx.c0.rspValid && isUmsgResponse(ccip_rx.c0.hdr.resp_type)) begin
	    if (C0RxUMsgHdr.umsg_type) begin
	       if (cfg.enable_cl_view) $display("%d\t   \tUMsgHint   \t%d\n",
						$time,
						C0RxUMsgHdr.umsg_id
						);
	       $fwrite(log_fd, "%d\t   \tUMsgHint   \t%d\n",
		       $time,
		       C0RxUMsgHdr.umsg_id
		       );
	    end
	    else if (~C0RxUMsgHdr.umsg_type) begin
	       if (cfg.enable_cl_view) $display("%d\t   \tUMsgData   \t%d\t%x\n",
						$time,
						C0RxUMsgHdr.umsg_id,
						ccip_rx.c0.data
						);
	       $fwrite(log_fd, "%d\t   \tUMsgData   \t%d\t%x\n",
		       $time,
		       C0RxUMsgHdr.umsg_id,
		       ccip_rx.c0.data
		       );
	    end
	 end
	 // /**************** MEM -> AFU Interrupt Response  **************/
	 // if (C0RxIntrValid) begin
	 // end
	 //////////////////////// C1 RX CHANNEL TRANSACTIONS //////////////////////////
	 /****************** MEM -> AFU Write Response  ****************/
	 if (ccip_rx.c1.rspValid && isWrLineResponse(ccip_rx.c1.hdr.resp_type)) begin
	    if (cfg.enable_cl_view) $display("%d\t%s\t%s\t%x\t%s",
	 				     $time,
	 				     print_channel(ccip_rx.c1.hdr.vc_used),
	 				     print_c1_resptype(ccip_rx.c1.hdr.resp_type),
	 				     ccip_rx.c1.hdr.mdata,
					     print_clnum(ccip_rx.c1.hdr.cl_num));
	    $fwrite(log_fd, "%d\t%s\t%s\t%x\t%s\n",
	 	    $time,
	 	    print_channel(ccip_rx.c1.hdr.vc_used),
	 	    print_c1_resptype(ccip_rx.c1.hdr.resp_type),
	 	    ccip_rx.c1.hdr.mdata,
		    print_clnum(ccip_rx.c1.hdr.cl_num));
	 end
	 if (ccip_rx.c1.rspValid && isWrFenceResponse(ccip_rx.c1.hdr.resp_type)) begin
	    if (cfg.enable_cl_view) $display("%d\t%s\tWrFenceRsp\t%x",
					     $time,
					     print_channel(ccip_rx.c1.hdr.vc_used),
					     ccip_rx.c1.hdr.mdata);
	    $fwrite(log_fd, "%d\t%s\tWrFenceRsp\t%x\n",
		    $time,
		    print_channel(ccip_rx.c1.hdr.vc_used),
		    ccip_rx.c1.hdr.mdata);
	 end
	 // /**************** MEM -> AFU Interrupt Response  **************/
	 // if (C1RxIntrValid) begin
	 // end
	 ////////////////////////////// FINISH command ////////////////////////////////
	 if (finish_logger == 1) begin
	    $fclose(log_fd);
	 end
	 //////////////////////////////////////////////////////////////////////////////
	 // Wait till next clock
	 $fflush(log_fd);
	 @(posedge clk);
      end
   end

endmodule
