mcadler@vs-fpga-5.hd.intel.com.75942:1450824863